rom(0) <= "11100011101000000000000000000000"
rom(1) <= 11100011101000000001000000000001
rom(2) <= 11100011101000000010000000000001
rom(3) <= 11100101100000000001000000000001
rom(4) <= 11100101100000000010000000000010
rom(5) <= 11100001101000000001000000000001
rom(6) <= 11100001101000000001000000000001
rom(7) <= 11100001101000000001000000000001
rom(8) <= 11100001101000000001000000000001
rom(9) <= 11100001101000000001000000000001
rom(10) <= 11100001101000000001000000000001
rom(11) <= 11100001101000000001000000000001
rom(12) <= 11100001101000000001000000000001
rom(13) <= 11100001101000000001000000000001
rom(14) <= 11100001101000000001000000000001
rom(15) <= 11100001101000000001000000000001
rom(16) <= 11100001101000000001000000000001
rom(17) <= 11100001101000000001000000000001
rom(18) <= 11100001101000000001000000000001
rom(19) <= 11100001101000000001000000000001
rom(20) <= 11100001101000000001000000000001
rom(21) <= 11100001101000000001000000000001
rom(22) <= 11100001101000000001000000000001
rom(23) <= 11100001101000000001000000000001
rom(24) <= 11100001101000000001000000000001
rom(25) <= 11100001101000000001000000000001
rom(26) <= 11100001101000000001000000000001
rom(27) <= 11100001101000000001000000000001
rom(28) <= 11100001101000000001000000000001
rom(29) <= 11100001101000000001000000000001
rom(30) <= 11100001101000000001000000000001
rom(31) <= 11100001101000000001000000000001
rom(32) <= 11100001101000000001000000000001
rom(33) <= 11100001101000000001000000000001
rom(34) <= 11100001101000000001000000000001
rom(35) <= 11100001101000000001000000000001
rom(36) <= 11100001101000000001000000000001
rom(37) <= 11100001101000000001000000000001
rom(38) <= 11100001101000000001000000000001
rom(39) <= 11100001101000000001000000000001
rom(40) <= 11100001101000000001000000000001
rom(41) <= 11100001101000000001000000000001
rom(42) <= 11100001101000000001000000000001
rom(43) <= 11100001101000000001000000000001
rom(44) <= 11100001101000000001000000000001
rom(45) <= 11100001101000000001000000000001
rom(46) <= 11100001101000000001000000000001
rom(47) <= 11100001101000000001000000000001
rom(48) <= 11100001101000000001000000000001
rom(49) <= 11100001101000000001000000000001
rom(50) <= 11100001101000000001000000000001
rom(51) <= 11101010111111111111111111010000
rom(52) <= 111010101111111111111111110100
