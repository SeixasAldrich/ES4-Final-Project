library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity progrom is

	port(
		addr : in unsigned(31 downto 0);
		data : out std_logic_vector(31 downto 0)
		);

end;

architecture synth of progrom is

begin



end;
